test
test
test this is a 
test
